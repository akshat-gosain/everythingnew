`include "full_adder.v"
module ripple_carry_4_bit_adder (input [3:0] A, input [3:0] B, input C0, output [3:0] Sum, output C4)



endmodule
