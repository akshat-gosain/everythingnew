module half_adder (input x, input y, output S, output C)



endmodule
