module D_ff(input clk, input reset, input D, output reg Q)



endmodule